module simplewire(
    input in, output out 
);

    assign out = in; // 출력 = 입력 

endmodule