module simplewire(
    input in,
    output out
);

    assign out = in;

endmodule
