module modulepos(

    input a, b, c, d, 
    output out1, out2

);

    mod_a ( out1, out2, a, b, c, d);

endmodule