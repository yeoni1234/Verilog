module modules(

input a, b,
output out

);


endmodule