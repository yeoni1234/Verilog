module modules(

input a, b,
output out

);

    mod_a (a, b, out);
    
    //mod_a ( .in1(a), .in2(b), .out(out));

endmodule

