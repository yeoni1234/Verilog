module top_module(zero);
    
    output zero;

endmodule