module alwayscase(

    input [2:0] sel, 
    input [3:0] data0,
    input [3:0] data1,
    input [3:0] data2,
    input [3:0] data3,
    input [3:0] data4,
    input [3:0] data5,
    output reg [3:0] out


);

    always @(*) begin

        case (sel)
            3'b000 : out = data0;
            3'b001 : out = data1;
            3'b010 : out = data2;
            3'b011 : out = data3;
            3'b100 : out = data4;
            3'b101 : out = data5;

            default : out = 0; // case 문을 사용할 때는 default값을 적어줌으로써 latch방지!
        endcase
    end
    

endmodule