module vectorgates(

    input [2:0] a, b,
    output [2:0] out_or_bitwise,
    output out_or_logical,
    output [5:0] out_not
);



endmodule