module moduleshift8(

    input clk,
    input [7:0] d,
    input [1:0] sel,
    output [7:0] q
);



endmodule