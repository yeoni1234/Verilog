module faad(

    input a, b, cin,
    output cout, sum

);

    always @(*) begin


    end

endmodule