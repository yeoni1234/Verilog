module abc( output one );


    assign one = 1; //1'b1;

endmodule

